magic
tech sky130A
magscale 1 2
timestamp 1716650568
<< pwell >>
rect 2924 244 4654 328
rect 8904 104 14430 172
rect 13206 102 14430 104
rect 8906 -314 9996 -244
rect 13996 -314 14428 102
rect 9564 -446 9996 -314
rect 9564 -512 14430 -446
rect 8908 -718 9998 -648
rect 13998 -718 14430 -512
rect 9566 -872 9998 -718
rect 13998 -872 14430 -868
rect 9564 -938 14430 -872
rect 8908 -1138 9998 -1068
rect 13998 -1138 14430 -938
rect 9566 -1280 9998 -1138
rect 13996 -1280 14428 -1278
rect 3020 -1378 4530 -1344
rect 9566 -1346 14428 -1280
rect 8906 -1544 9996 -1474
rect 13996 -1544 14428 -1346
rect 9564 -1688 9996 -1544
rect 9564 -1754 14426 -1688
rect 8904 -1958 9994 -1888
rect 13994 -1958 14426 -1754
rect 9562 -2088 9994 -1958
rect 9562 -2154 14424 -2088
rect 8902 -2354 9992 -2284
rect 13992 -2354 14424 -2154
rect 9560 -2540 9992 -2354
rect 8906 -2746 9996 -2676
rect 13996 -2746 14428 -2490
rect 4578 -3224 5840 -3222
rect 4578 -3226 8204 -3224
rect 14492 -3226 14594 -78
rect 4578 -3270 14594 -3226
rect 2924 -3286 14594 -3270
rect 2924 -3288 5840 -3286
rect 10536 -3288 14594 -3286
<< viali >>
rect 3020 268 4530 302
rect 3020 -28 4530 6
rect 3020 -148 4530 -114
rect 14524 -348 14558 -210
rect 3020 -444 4530 -410
rect 3020 -552 4530 -518
rect 14526 -752 14560 -614
rect 3020 -848 4530 -814
rect 3020 -972 4530 -938
rect 14526 -1172 14560 -1034
rect 3020 -1268 4530 -1234
rect 3020 -1378 4530 -1344
rect 14524 -1578 14558 -1440
rect 3020 -1674 4530 -1640
rect 3020 -1792 4530 -1758
rect 14522 -1992 14556 -1854
rect 3020 -2088 4530 -2054
rect 3020 -2188 4530 -2154
rect 14520 -2388 14554 -2250
rect 3020 -2484 4530 -2450
rect 3020 -2580 4530 -2546
rect 14524 -2780 14558 -2642
rect 3020 -2876 4530 -2842
rect 3020 -2976 4530 -2942
rect 3020 -3272 4530 -3238
<< metal1 >>
rect 2924 302 4654 328
rect 2924 268 3020 302
rect 4530 268 4654 302
rect 2924 244 4654 268
rect 6 38 904 238
rect 184 36 904 38
rect 2924 6 4652 244
rect 8904 104 14430 172
rect 13206 102 14430 104
rect 2924 -28 3020 6
rect 4530 -28 4652 6
rect 2924 -114 4652 -28
rect 2924 -148 3020 -114
rect 4530 -148 4652 -114
rect 6 -390 906 -190
rect 2924 -410 4652 -148
rect 13996 -28 14430 102
rect 8906 -314 9996 -244
rect 13996 -314 14428 -28
rect 14492 -210 14594 -78
rect 2924 -444 3020 -410
rect 4530 -444 4652 -410
rect 2924 -518 4652 -444
rect 9564 -446 9996 -314
rect 14492 -348 14524 -210
rect 14558 -348 14594 -210
rect 9564 -512 14430 -446
rect 2924 -552 3020 -518
rect 4530 -552 4652 -518
rect 6 -786 908 -586
rect 2924 -814 4652 -552
rect 8908 -718 9998 -648
rect 13998 -718 14430 -512
rect 14492 -614 14594 -348
rect 2924 -848 3020 -814
rect 4530 -848 4652 -814
rect 2924 -938 4652 -848
rect 9566 -872 9998 -718
rect 14492 -752 14526 -614
rect 14560 -752 14594 -614
rect 13998 -872 14430 -868
rect 9564 -938 14430 -872
rect 2924 -972 3020 -938
rect 4530 -972 4652 -938
rect 6 -1208 908 -1008
rect 2924 -1234 4652 -972
rect 8908 -1138 9998 -1068
rect 13998 -1138 14430 -938
rect 14492 -1034 14594 -752
rect 2924 -1268 3020 -1234
rect 4530 -1268 4652 -1234
rect 2924 -1344 4652 -1268
rect 2924 -1378 3020 -1344
rect 4530 -1378 4652 -1344
rect 9566 -1280 9998 -1138
rect 14492 -1172 14526 -1034
rect 14560 -1172 14594 -1034
rect 13996 -1280 14428 -1278
rect 9566 -1346 14428 -1280
rect 6 -1592 906 -1392
rect 2924 -1640 4652 -1378
rect 8906 -1544 9996 -1474
rect 13996 -1544 14428 -1346
rect 14492 -1440 14594 -1172
rect 2924 -1674 3020 -1640
rect 4530 -1674 4652 -1640
rect 2924 -1758 4652 -1674
rect 9564 -1688 9996 -1544
rect 14492 -1578 14524 -1440
rect 14558 -1578 14594 -1440
rect 9564 -1754 14426 -1688
rect 2924 -1792 3020 -1758
rect 4530 -1792 4652 -1758
rect 6 -2026 904 -1826
rect 2924 -2054 4652 -1792
rect 8904 -1958 9994 -1888
rect 13994 -1958 14426 -1754
rect 14492 -1854 14594 -1578
rect 2924 -2088 3020 -2054
rect 4530 -2088 4652 -2054
rect 2924 -2154 4652 -2088
rect 9562 -2088 9994 -1958
rect 14492 -1992 14522 -1854
rect 14556 -1992 14594 -1854
rect 9562 -2154 14424 -2088
rect 2924 -2188 3020 -2154
rect 4530 -2188 4652 -2154
rect 0 -2406 902 -2206
rect 2924 -2450 4652 -2188
rect 8902 -2354 9992 -2284
rect 13992 -2354 14424 -2154
rect 14492 -2250 14594 -1992
rect 2924 -2484 3020 -2450
rect 4530 -2484 4652 -2450
rect 2924 -2546 4652 -2484
rect 9560 -2490 9992 -2354
rect 14492 -2388 14520 -2250
rect 14554 -2388 14594 -2250
rect 9560 -2540 14428 -2490
rect 2924 -2580 3020 -2546
rect 4530 -2580 4652 -2546
rect 0 -2814 906 -2614
rect 2924 -2842 4652 -2580
rect 2924 -2876 3020 -2842
rect 4530 -2876 4652 -2842
rect 2924 -2942 4652 -2876
rect 2924 -2976 3020 -2942
rect 4530 -2976 4652 -2942
rect 2924 -3000 4652 -2976
rect 0 -3200 4652 -3000
rect 8906 -2746 9996 -2676
rect 13996 -2746 14428 -2540
rect 14492 -2642 14594 -2388
rect 8906 -3142 9334 -2746
rect 14492 -2780 14524 -2642
rect 14558 -2780 14594 -2642
rect 842 -3202 4652 -3200
rect 2924 -3222 4652 -3202
rect 2924 -3224 5840 -3222
rect 2924 -3226 8204 -3224
rect 14492 -3226 14594 -2780
rect 2924 -3238 14594 -3226
rect 2924 -3272 3020 -3238
rect 4530 -3272 14594 -3238
rect 2924 -3286 14594 -3272
rect 2924 -3288 5840 -3286
rect 10536 -3288 14594 -3286
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR1
timestamp 1716578501
transform 0 1 4902 -1 0 -3107
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR2
timestamp 1716578501
transform 0 1 4906 -1 0 -279
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR3
timestamp 1716578501
transform 0 1 4908 -1 0 -683
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR4
timestamp 1716578501
transform 0 1 4908 -1 0 -1103
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR5
timestamp 1716578501
transform 0 1 4906 -1 0 -1509
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR6
timestamp 1716578501
transform 0 1 4904 -1 0 -1923
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR7
timestamp 1716578501
transform 0 1 4902 -1 0 -2319
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR8
timestamp 1716578501
transform 0 1 4906 -1 0 -2711
box -201 -4598 201 4598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR9
timestamp 1716578501
transform 0 1 11996 -1 0 -279
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR10
timestamp 1716578501
transform 0 1 11998 -1 0 -683
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR11
timestamp 1716578501
transform 0 1 11998 -1 0 -1103
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR12
timestamp 1716578501
transform 0 1 11996 -1 0 -1509
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR13
timestamp 1716578501
transform 0 1 11994 -1 0 -1923
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR14
timestamp 1716578501
transform 0 1 11992 -1 0 -2319
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR15
timestamp 1716578501
transform 0 1 11996 1 0 -2711
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_3KK54B  XR16
timestamp 1716578501
transform 0 1 4904 -1 0 137
box -201 -4598 201 4598
<< labels >>
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 GND
port 8 nsew
flabel metal1 0 -2814 200 -2614 0 FreeSans 256 0 0 0 b0
port 0 nsew
flabel metal1 0 -2406 200 -2206 0 FreeSans 256 0 0 0 b1
port 1 nsew
flabel metal1 6 -2026 206 -1826 0 FreeSans 256 0 0 0 b2
port 2 nsew
flabel metal1 6 -1592 206 -1392 0 FreeSans 256 0 0 0 b3
port 3 nsew
flabel metal1 6 -1208 206 -1008 0 FreeSans 256 0 0 0 b4
port 4 nsew
flabel metal1 6 -786 206 -586 0 FreeSans 256 0 0 0 b5
port 5 nsew
flabel metal1 6 -390 206 -190 0 FreeSans 256 0 0 0 b6
port 6 nsew
flabel metal1 6 38 206 238 0 FreeSans 256 0 0 0 b7
port 7 nsew
flabel metal1 14230 -28 14430 172 0 FreeSans 256 0 0 0 OUT
port 9 nsew
<< end >>
